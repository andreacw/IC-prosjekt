[aimspice]
[description]
1720
Analog circuit PROJECT(1 pixel)

.param Wn={2u} 
.param Wp={2u}
.param Ln={0.7u}
.param Lp={0.7u}
.param Cs={0.6pf}
.param cc1={3pf}
.param T= 10m
.param PW = {T/2}
.param TRF = {T/100}
.param Ipd_1 = 200p

V_EXP gEXPOSE 0 dc PULSE(1.8 0 5m TRF TRF PW T)
V_ERASE gERASE 0 dc PULSE(1.8 0 10m TRF TRF PW T)
V_NRE gNRE 0 dc PULSE(0 0 15m TRF TRF PW T)
VDD vdd 0 dc 1.8v
*-------------------------------------------------------
*.plot tran(gEXPOSE) v(gERASE) v(N2)
.plot tran(gNRE) v(OUT) v(N2) V(gEXPOSE)

*X2 gEXPOSE gERASE vdd N2 del_1
*X3 N2 gNRE vdd OUT del_2
X1 vdd gExpose gErase gNRE OUT N2 onePixel
X4 vdd OUT del_3 

*------------------------------------------------------
.subckt  del_1 gEXPOSE gERASE vdd N2
X1 vdd N1 PhotoDiode
MN1 N1 gEXPOSE N2 0 NMOS L=Ln W=Wn
MN2 N2 gERASE 0 0 NMOS L=Ln W=Wn
CS N2 0 Cs
.ends 

*------------------------------------------------------
.subckt del_2 N2 gNRE vdd OUT1
MP3 0 N2 N3 vdd PMOS L=Lp W=Wp
MP4 N3 gNRE OUT1 vdd PMOS L=Lp W=Wp
.ends

*------------------------------------------------------
.subckt onePixel vdd gExpose gErase gNRE N2 OUT1
	X2 gEXPOSE gERASE vdd N2 del_1
	X3 N2 gNRE vdd OUT1 del_2
.ends

*------------------------------------------------------
.subckt del_3 vdd OUT1
MP5 OUT1 OUT1 vdd vdd PMOS W=Wp L=Lp
CC1 OUT1 0 cc1
.ends 

*------------------------------------------------------
.subckt PhotoDiode  VDD N1_R1C1 
I1_R1C1  VDD   N1_R1C1   DC  Ipd_1
d1 N1_R1C1 vdd dwell 1
.model dwell d cj0=1e-14 is=1e-12 m=0.5 bv=40
Cd1 N1_R1C1 VDD 30f
.ends 


.include C:\Users\haral\OneDrive\NTNU\IC\Project\p18_cmos_models_tt.inc
.include C:\Users\haral\OneDrive\NTNU\IC\Project\p18_model_card.inc

[tran]
0.1m
50m
X
X
0
[ana]
4 0
[end]
