[aimspice]
[description]
544
Analog part , IC prosjekt

.include p18_cmos_models.inc
.include p18_model_card.inc

VDD vdd 0 dc 1.8V

.param EXPOSE = 0.5s
.param EREASE = 0
.param MP1W = 2.6u
.param MP1L = 0.6u

* Photo diode
.subckt PhotoDiode  VDD N1_R1C1 
I1_R1C1  VDD   N1_R1C1   DC  Ipd_1
d1 N1_R1C1 vdd dwell 1
.model dwell d cj0=1e-14 is=1e-12 m=0.5 bv=40
Cd1 N1_R1C1 VDD 30f
.ends

* MN1 DRAIN GATE SOURCE BULK NMOS WIDTH LENGTH 
* MP1 SOURCE GATE DRAIN BULK PMOS WIDTH LENGTH

PD1 PhotoDiode VDD N1
MP1 N2 EXPOSE N1 VSS PMOS MP1W MP1L 



[end]
